module DE1_SoC ();
endmodule
